module mips(
    input logic clk, reset, addr, mem_write,
    input logic [31:0] read_data,

    output logic [31:0] write_data
);

    

endmodule