module main_decoder();


endmodule