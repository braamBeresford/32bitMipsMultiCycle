module alu_decoder();


endmodule